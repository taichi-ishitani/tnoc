`ifndef NOC_BFM_STATUS_SVH
`define NOC_BFM_STATUS_SVH
typedef tue_status_dummy  noc_bfm_status;
`endif
