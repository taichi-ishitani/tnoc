`ifndef TNOC_BFM_PKG_SV
`define TNOC_BFM_PKG_SV
package tnoc_bfm_pkg;
  import  uvm_pkg::*;
  import  tue_pkg::*;
  import  tnoc_bfm_types_pkg::*;

  `include  "uvm_macros.svh"
  `include  "tue_macros.svh"
  `include  "tnoc_bfm_macro.svh"

  typedef virtual tnoc_bfm_flit_if  tnoc_bfm_flit_vif;

  `include  "tnoc_bfm_configuration.svh"
  `include  "tnoc_bfm_status.svh"
  `include  "tnoc_bfm_flit_item.svh"
  `include  "tnoc_bfm_packet_item.svh"

  `include  "tnoc_bfm_component_base.svh"
  `include  "tnoc_bfm_packet_monitor.svh"
  `include  "tnoc_bfm_packet_sequencer.svh"
  `include  "tnoc_bfm_packet_driver.svh"
  `include  "tnoc_bfm_packet_agent.svh"
endpackage
`endif
