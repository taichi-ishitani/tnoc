import  tnoc_config_pkg::*,
        tnoc_enums_pkg::tnoc_port_type,
        tnoc_enums_pkg::TNOC_LOCAL_PORT,
        tnoc_enums_pkg::TNOC_INTERNAL_PORT,
        tnoc_enums_pkg::is_local_port,
        tnoc_enums_pkg::is_internal_port;
