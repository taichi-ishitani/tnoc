`ifndef TNOC_CONFIG_DEFINES_SVH
`define TNOC_CONFIG_DEFINES_SVH

`ifndef TNOC_DEFAULT_ADDRESS_WIDTH
  `define TNOC_DEFAULT_ADDRESS_WIDTH  64
`endif

`ifndef TNOC_MAX_DATA_WIDTH
  `define TNOC_MAX_DATA_WIDTH 256
`endif

`ifndef TNOC_DEFAULT_DATA_WIDTH
  `define TNOC_DEFAULT_DATA_WIDTH `TNOC_MAX_DATA_WIDTH
`endif

`ifndef TNOC_DEFAULT_ID_X_WIDTH
  `define TNOC_DEFAULT_ID_X_WIDTH 5
`endif

`ifndef TNOC_DEFAULT_ID_Y_WIDTH
  `define TNOC_DEFAULT_ID_Y_WIDTH 5
`endif

`ifndef TNOC_DEFAULT_VIRTUAL_CHANNELS
  `define TNOC_DEFAULT_VIRTUAL_CHANNELS 2
`endif

`ifndef TNOC_DEFAULT_TAGS
  `define TNOC_DEFAULT_TAGS 256
`endif

`ifndef TNOC_DEFAULT_MAX_BURST_LENGTH
  `define TNOC_DEFAULT_MAX_BURST_LENGTH 256
`endif

`ifndef TNOC_DEFAULT_FIFO_DEPTH
  `define TNOC_DEFAULT_FIFO_DEPTH 8
`endif

`ifndef TNOC_DEFAULT_SIZE_X
  `define TNOC_DEFAULT_SIZE_X 3
`endif

`ifndef TNOC_DEFAULT_SIZE_Y
  `define TNOC_DEFAULT_SIZE_Y 3
`endif

`ifndef TNOC_DEFAULT_ERROR_DATA
  `define TNOC_DEFAULT_ERROR_DATA '1
`endif

`endif
