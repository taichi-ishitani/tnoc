`ifndef NOC_BFM_MACROS_SVH
`define NOC_BFM_MACROS_SVH

`ifndef NOC_BFM_MAX_ADDRESS_WIDTH
  `define NOC_BFM_MAX_ADDRESS_WIDTH 64
 `endif

`ifndef NOC_BFM_MAX_DATA_WIDTH
  `define NOC_BFM_MAX_DATA_WIDTH  256
`endif

`ifndef NOC_BFM_MAX_ID_X_WIDTH
  `define NOC_BFM_MAX_ID_X_WIDTH  8
`endif

`ifndef NOC_BFM_MAX_ID_Y_WIDTH
  `define NOC_BFM_MAX_ID_Y_WIDTH  8
`endif

`ifndef NOC_BFM_MAX_TAG_WIDTH
  `define NOC_BFM_MAX_TAG_WIDTH 8
`endif

`ifndef NOC_BFM_MAX_LENGTH_WIDTH
  `define NOC_BFM_MAX_LENGTH_WIDTH  5
`endif

`endif
