import  tnoc_config_pkg::*,
        tnoc_enums_pkg::*;
